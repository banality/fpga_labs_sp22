`timescale 1ns/1ns
`include "adder.vh"

`define SECOND 1000000000
`define MS 1000000

module adder_testbench();
    reg [`ADDER_BIT_WIDTH-1:0] a;
    reg [`ADDER_BIT_WIDTH-1:0] b;
    wire [`ADDER_BIT_WIDTH:0] sum;

    structural_adder sa (
        .a(a),
        .b(b),
        .sum(sum)
    );

    integer ai, bi;
    initial begin
        `ifdef IVERILOG
            $dumpfile("adder_testbench.fst");
            $dumpvars(0, adder_testbench);
        `endif
        `ifndef IVERILOG
            $vcdpluson;
        `endif

        // for (ai = 0; ai <=10024; ai = ai+1) begin
        //     for (bi = 0; bi <=10024; bi = bi+1) begin
        //         a = ai;
        //         b = bi;
        //         #(2);
        //     end
        // end

        a = $urandom();
        b = $urandom();
        #(2);

        a = 14'd1;
        b = 14'd1;
        #(2);
        if (sum != 15'd2) $display("ERROR: Expected sum to be 2, actual value: %d", sum);

        a = 14'd0;
        b = 14'd1;
        #(2);
        if(sum != 15'd1) $display("ERROR: Expected sum to be 1, actual value: %d", sum);

        a = 14'd10;
        b = 14'd10;
        #(2);
        if (sum != 15'd20) begin
            $error("Expected sum to be 20, a: %d, b: %d, actual value: %d", a, b, sum);
            $fatal(1);
        end

        `ifndef IVERILOG
            $vcdplusoff;
        `endif
        $finish();
    end
endmodule
