`define ADDER_BIT_WIDTH 32
